`ifndef DEFS_DONE
`define DEFS_DONE
package defs;
	parameter CPUID   = "SI MIPS YO";
	parameter VERSION = "0.9       ";

endpackage

import defs::*;

`endif